----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:00:16 08/21/2014 
-- Design Name: 
-- Module Name:    bitadder - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity bitadder is
    Port ( A : in  STD_LOGIC;
           B : in  STD_LOGIC;
			  Cin : in STD_LOGIC;
           Cout : out  STD_LOGIC;
           S : out  STD_LOGIC);
end bitadder;

architecture Behavioral of bitadder is

begin

	S <= A xor B xor Cin;
	Cout <= (A and B) or (Cin and (A xor B));

end Behavioral;

